----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Fernando Leon
-- 
-- Create Date:    15:02:45 03/20/2024 
-- Design Name: 
-- Module Name:    toggler - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity toggler is
    Port ( t : in  STD_LOGIC;
           o : out  STD_LOGIC);
end toggler;

architecture Behavioral of toggler is
	signal s: STD_LOGIC := '0';
begin
	process(t,s)
	begin
		if rising_edge(t) then
			s <= not s;
		end if;
		o <= s;
	end process;


end Behavioral;

